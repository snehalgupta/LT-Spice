*Question4
V1 1 0 AC 1
R1 2 1 0.0796k
R2 3 2 0.0796k
C1 4 2 1u
e 4 0 3 5 999k
C2 0 3 1u
R3 5 4 10k
R4 0 5 5.55k
R5 0 4 10k
.ac dec 100 1 10k
.end