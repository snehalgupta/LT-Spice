* Question 3
V1 1 0 80;
R1 1 2 20;
R2 0 2 20;
L1 2 0 15 ic=0;
C1 2 0 0.0333 ic=0;

.op
.tran 0.001 10 uic
.end
