* question2
r1 0 1 4k
r2 1 2 12k
c1 3 4 0.047u
r3 4 5 1k
r4 2 5 11.11k
vi 3 5 AC 1
e 2 0 1 4 999k
.ac dec 100 1 100k
.ends

