* Question 4
L1 0 1 2 ic=3;
R1 0 1 8;
C1 1 0 0.25 ic=24;
.op
.tran 0.01 50 uic
.end
