* question1
v1 1 0 sin(0 40 1 0 0 0 1)
r1 1 2 8
c1 1 2 0.5
l1 2 3 4
v2 3 0 sin(0 20 0.159 0 90 0 1)
.tran 1 100
