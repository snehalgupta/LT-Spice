//if
V1 1 0 pwl(0 24 0.01 0)
R1 1 2 4
R2 2 0 4
l3 2 3 4
R4 3 0 8
.tran 1 10
.end