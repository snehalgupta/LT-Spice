*Q2
V1 1 0 AC 100.
R1  1 2 1000
C1 2 0 1m
R2 2 3 1000
G1 3 0 2 0 0.1
R3 3 4 1000
L1 4 0 1m

.ac dec 100 1 10k
.end