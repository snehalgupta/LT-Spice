* Question 2
V1 1 0 80
R1 1 2 160
R2 2 3 80
H1 3 0 V1 80
V2 2 4 PWL(0 80 0.01m 0)
L1 4 0 30
R3 4 0 40
C1 4 0 0.01666
.tran 14
.end
