* question1
r1 0 1 10k
r2 1 3 10k
r3 2 0 1k
c1 2 4 1u
vi 4 0 AC 1
e 3 0 1 2 999k
.ac dec 100 1 100k
.ends

