* circuit2
R1 1 0 5
V1 2 1 8V
R2 2 0 2
V2 3 2 4V
R3 2 4 4
R4 3 0 4
R5 3 4 1
V3 4 0 10V
.op
.end 
