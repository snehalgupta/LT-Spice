*Question3
R1 1 0 25k
R2 4 1 20k
e 4 0 1 3 999k
C1 3 0 0 0.047u
V1 6 0 AC 1
R3 3 5 1.54k
C2 5 4 0.047u
R4 5 6 1.54k
R5 4 0 10k
.ac dec 100 1 10k
.end

