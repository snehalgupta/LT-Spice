* Question 4
V1 1 0 10V;
C1 1 2 47u ic=0;
C2 1 2 20u ic=0;
R1 2 0 3k;

.op
.tran 0.05 1 uic
.end